location Nice is "Port de Villefranche-sur-Mer, France"
location Cerbre is "Cape Cerbre France"
location Toulon is "Toulon France"
location Hyeres is "Hyeres France"
location Frejus is "Frejus France"
location Antibes is "Antibes France"
location Cannes is "Cannes France"
location Vendres is "Port Vendres"
location Monaco is "Monaco"
