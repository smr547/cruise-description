vessel Trilogy name: "Trilogy" flag: "Australia" rego: 12345

location Sant_Carles is "Sant Carles de la Rapita"
location Barcelona is "Port of Barcelona Spain"
location Blanes is "Blanes Spain"
location WPa at 6.7 43.2 is "a waypoint"
location Roses is "Roses Spain"
location Menton is "Menton Italy"
location Cerbre is "Cape Cerbre France"
location Vendres is "Port Vendres"
location Bastia is "Bastia Corsica"
location Calvi is "Calvi Corsica"
location Macinaggio is "Macinaggio Corsica"
location Propriano is "Propriano Corsica"
location Banifacio is "Banifacio Corsica"
location Porto_Vecchio is "Porto Vecchio Corsica"
location ST_FLOR is "St Florent Corsica"
location Alghero is "Alghero Sardinia"
location Arbatax is "Arbatax Sardinia"
location Cagliari is "Cagliari Sardinia"
location Calsetta is "Calasetta Sardinia"
location Carloforte is "Carloforte Sardinia"
location Castelsardo is "Castelsardo Sardina"
location Rossa is "Isola Rossa Sardina"
location Maddalena is "Maddalena Archipelago Sardina"
location Olbia is "Olbia Sardinia"
location Cervo is "Porto Cervo Sardinia"
location Torres is "Porto Torres Sardinia"
location Portoscuso is "Portoscuso Sardinia"
location Gallura is "Santa Teresa Gallura Sardinia"
location Torregrande is "Torregrande  Sardinia"
location Tuelada is "Tuelada Sardinia"
location Villasimius is "Villasimius Sardinia"
location La_Spezia is "La Spezia Italy"
location Termini is "Termini Italy"
location Fanciullo is "Fanciullo Italy"

person smr name: "Steven Michael Ring"
person isf name: "Irene Sarrah Farthing"

season Steven_cruise vessel Trilogy

cruise  "Shakedown"
	Sant_Carles
        crew smr joins on 31/3/19 as skipper
        crew wp  joins on 07/4/19 as mate
	Tarragona for 1 night
	Barcelona for 4 nights
        crew wp leaves
cruise  "Barcelona to Nice"
	Barcelona
	Blanes
	Roses
	Cerbre
	Vendres
	Toulon
	Hyeres
	WPa
	Frejus
	Cannes
	Nice
cruise  "Nice to Naples via Corsica and Sardinia"
	Nice
	Monaco
	Menton
	Imperia
	Calvi
	Propriano
	Banifacio
	Gallura
	Maddalena
	Cervo
	Arbatax
	Cagliari
	Capri
	Naples
cruise  "Naples to Genoa via Amalfi Coast and Cinque Terre"
	Naples
	Sorrento
	Termini
	Amalfi
	Salerno
	Capri
	Ischia
	Formia
	Anzio
	Ostia
	Fanciullo
	Orbetello
	Follonica
	Piombino
	Portoferraio
	Livorno
	La_Spezia
	Chiavari
	Genoa
