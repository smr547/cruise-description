vessel Trilogy name: "Trilogy" flag: "Australia" rego: 12345 speed: 7.5

location WPa at 6.7 43.2 is "a waypoint"
location WPb at 6.7 43.3 is "a waypoint"

use https://smr547.github.io/locations/corsica.txt
use https://smr547.github.io/locations/france_med_coast.txt
use https://smr547.github.io/locations/sardinia.txt
use https://smr547.github.io/locations/italy.txt
use https://smr547.github.io/locations/spain_med_coast.txt

use file:///home/smring/projects/cruise-description/grammar/people.cdl


season Steven_cruise vessel Trilogy begins in Sant_Carles

cruise  "Shakedown" departs Sant_Carles on 14/4/19 at 1000
	Sant_Carles
        crew smr joins on 31/3/19 as skipper in Sant_Carles
        crew wp  joins on 08/4/19 as mate in Sant_Carles
	Tarragona for 1 night
	Barcelona for 4 nights
        crew wp leaves on 16/4/19

cruise  "Barcelona to Nice" departs Barcelona on 17/4/19 at 1000
        crew gh joins on 16/4/19 in Barcelona
        crew cm joins on 16/4/19 in Barcelona
        crew sjr joins on 16/4/19 in Barcelona
        crew pjr joins on 16/4/19 in Barcelona
        crew ar joins on 16/4/19 in Barcelona
	Barcelona
	Blanes for 1 night
	Roses for 2 night
	Cerbre for 1 night
	Vendres for 2 night
	Toulon for 1 night
	Hyeres for 1 night
	via WPa, WPb
	Frejus for 1 night
	Cannes for 1 night
        Antibes for 2 nights
	Nice for 4 nights
	crew gh leaves on 30/4/19 in Nice
	crew cm leaves on 30/4/19 in Nice
	crew sjr leaves on 1/5/19 in Nice
	crew ar leaves on 1/5/19 in Nice
	crew pjr leaves on 1/5/19 in Nice

cruise  "Nice to Naples via Corsica and Sardinia" departs Nice on 3/5/19 at 1000
	crew po joins on 1/5/19 as mate in Nice
	crew wp joins on 1/5/19 in Nice
	crew rb joins on 1/5/19 in Nice
	crew isf joins on 2/5/19 in Nice 
	Nice
	Monaco for 1 night
	Menton for 1 night
	Imperia for 1 night
	Calvi for 1 night
	Propriano for 1 night
	Banifacio for 1 night
	Gallura for 1 night
	Maddalena for 1 night
	Cervo for 1 night
	Arbatax for 1 night
	Cagliari for 1 night
	Capri for 1 night
	Naples for 1 night
	crew wp leaves on 2/6/19 in Naples
	crew rb leaves on 2/6/19 in Naples


cruise  "Naples to Genoa via Amalfi Coast and Cinque Terre" departs Naples on 4/6/19 at 1000
	crew kmt joins on 2/6/19 in Naples
	crew sgr joins on 2/6/19 in Naples
	Naples
	Sorrento for 1 night
	Termini for 1 night
	Amalfi for 1 night
	Salerno for 1 night
	Capri for 1 night
	Ischia for 1 night
	Formia for 1 night
	Anzio for 1 night
	Ostia for 1 night
	Fanciullo for 1 night
	Orbetello for 1 night
	Follonica for 1 night
	Piombino for 1 night
	Portoferraio for 1 night
	Livorno for 1 night
	La_Spezia for 1 night
	Chiavari for 1 night
	Genoa
	crew smr leaves on 30/6/19 in Genoa
	crew isf leaves on 30/6/19 in Genoa
	crew po leaves on 30/6/19 in Genoa
	crew kmt leaves on 30/6/19 in Genoa
	crew sgr leaves on 30/6/19 in Genoa
