vessel Trilogy name: "Trilogy" flag: "Australia" rego: 12345 speed: 7.5

#use http://ws.planacruise.online:5000/locations/corsica.txt
#use http://ws.planacruise.online:5000/locations/france_med_coast.txt
#use http://ws.planacruise.online:5000/locations/sardinia.txt
#use http://ws.planacruise.online:5000/locations/italy.txt
#use http://ws.planacruise.online:5000/locations/spain_med_coast.txt

use file:///Users/stevenring/projects/locations/docs/corsica.txt
use file:///Users/stevenring/projects/locations/docs/france_med_coast.txt
use file:///Users/stevenring/projects/locations/docs/sardinia.txt
use file:///Users/stevenring/projects/locations/docs/italy.txt
use file:///Users/stevenring/projects/locations/docs/spain_med_coast.txt
location Porquerolles is "Marina Porquerolles, France"
location Positano is "Positano, Italy"
location Portovenere is "Portovenere, Italy"
location Paraggi is "Paraggi, Italy"
location Cadaques is "Cadaques, Spain"
use file:///Users/stevenring/projects/cruise-description/grammar/people.cdl

season Steven_cruise vessel Trilogy begins in Sant_Carles

cruise  "Sant Carles to Nice" departs Sant_Carles on 2/5/19 at 1000
	Sant_Carles
        crew smr joins on 26/4/19 as skipper in Sant_Carles
        crew isf joins on 26/4/19 in Sant_Carles
        crew po  joins on 1/5/19 as mate in Sant_Carles
        Tarragona
        via Barcelona
        Blanes for 1 night
        Roses
        Cadaques for 1 night 
        Vendres for 1 nights
	Toulon for 1 night
	Porquerolles for 1 night
	Frejus for 1 night
        Antibes for 1 nights

cruise  "Antibes to Calvi" departs Antibes on 10/5/19 at 1000
	Antibes
	Calvi for 2 night

cruise  "Calvi to Sorrento via Corsica and Sardinia" departs Calvi on 16/5/19 at 1000
        Calvi
	crew wp joins on 15/5/19 in Calvi
	crew rb joins on 15/5/19 in Calvi
        via VI_2
        Crovani
        via Elbo, VI_3
        Girolata for 2 nights
        via Arone
        Cargese for 1 night
        via VI_4
        Ajaccio
        via VI_5
	Propriano for 2 night
        via VI_6, VI_7, VI_8
	Banifacio for 1 night
	Gallura for 1 night
	Maddalena for 1 night
	Cervo for 1 night
        Olbia for 1 night
	Capri for 1 night
	Sorrento for 1 night
	crew wp leaves on 2/6/19 in Sorrento
	crew rb leaves on 2/6/19 in Sorrento


cruise  "Sorrento to Genoa via Amalfi Coast and Cinque Terre" departs Sorrento on 4/6/19 at 1000
	crew kmt joins on 2/6/19 in Sorrento
	crew sgr joins on 2/6/19 in Sorrento
	Sorrento
        via IWP3_13, Positano
	Amalfi for 2 night
	Salerno for 1 night
	Capri for 1 night
	Ischia for 2 night
	Formia for 1 night
	Anzio for 1 night
	Fanciullo for 1 night
	Orbetello for 1 night
	Follonica for 1 night
	Piombino for 1 night
	Portoferraio for 2 night
	Livorno for 2 night
	La_Spezia for 1 night
        crew eif joins on 21/6/19 in La_Spezia
        via Portovenere
        Moneglia for 1 night
	Chiavari for 1 night
	Paraggi for 1 night
        Portofino for 2 nights
	Genoa
	crew smr leaves on 30/6/19 in Genoa
	crew isf leaves on 30/6/19 in Genoa
	crew po leaves on 30/6/19 in Genoa
	crew kmt leaves on 30/6/19 in Genoa
	crew sgr leaves on 30/6/19 in Genoa
	crew eif leaves on 30/6/19 in Genoa
