location Sant_Carles is Sant Carles de la Rapita
location Barcelona is Port of Barcelona Spain
location Blanes is Blanes Spain
location WPa at 6.7 43.2 is a waypoint
location Roses is Roses Spain
location Menton is Menton Italy
location Cerbre is Cape Cerbre France
location Vendres is Port Vendres

cruise (Shakedown 2019)
	Sant_Carles
	Tarragona
	Barcelona
	Blanes
	Roses
	Cerbre
	Vendres
	Toulon
	Hyeres
	WPa
	Frejus
	Cannes
	Nice
	Monaco
	Menton
	Imperia
	Calvi
