/Users/stevenring/projects/Trilogy/seasonal_plans/steven/steven_2020.cdl