location Sant_Carles is Sant Carles de la Rapita

cruise (Steven 2019)
	Sant_Carles
	Tarragona
	Barcelona
