location Sant_Carles is Sant Carles de la Rapita
location Tarragona is Tarragona, Spain
location Barcelona is Barcelona
