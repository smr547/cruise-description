location Sant_Carles is Sant Carles de la Rapita

cruise (Shakedown 2019)
	Sant_Carles
	Tarragona
	Barcelona
