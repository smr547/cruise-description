location Alghero is "Alghero Sardinia"
location Arbatax is "Arbatax Sardinia"
location Cagliari is "Cagliari Sardinia"
location Calsetta is "Calasetta Sardinia"
location Carloforte is "Carloforte Sardinia"
location Castelsardo is "Castelsardo Sardina"
location Rossa is "Isola Rossa Sardina"
location Maddalena is "Maddalena Archipelago Sardina"
location Olbia is "Olbia Sardinia"
location Cervo is "Porto Cervo Sardinia"
location Torres is "Porto Torres Sardinia"
location Portoscuso is "Portoscuso Sardinia"
location Gallura is "Santa Teresa Gallura Sardinia"
location Torregrande is "Torregrande  Sardinia"
location Tuelada is "Tuelada Sardinia"
location Villasimius is "Villasimius Sardinia"
