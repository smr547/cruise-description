vessel Trilogy name: "Trilogy" flag: "Australia" rego: 12345 speed: 7.5

use https://smr547.github.io/locations/corsica.txt
use https://smr547.github.io/locations/france_med_coast.txt
use https://smr547.github.io/locations/sardinia.txt
use https://smr547.github.io/locations/italy.txt
use https://smr547.github.io/locations/spain_med_coast.txt

use file:///Users/stevenring/projects/cruise-description/grammar/people.cdl

season Steven_cruise vessel Trilogy begins in Sant_Carles

cruise  "Sant Cales to Nice" departs Sant_Carles on 2/5/19 at 1000
	Sant_Carles
        crew smr joins on 30/4/19 as skipper in Sant_Carles
        crew isf joins on 30/4/19 as skipper in Sant_Carles
        crew po  joins on 1/4/19 as mate in Sant_Carles
	Toulon for 1 night
	Hyeres for 1 night
	Frejus for 1 night
        Antibes for 1 nights
	Cannes for 1 night
	Nice for 2 nights

cruise  "Nice to Naples via Corsica and Sardinia" departs Nice on 10/5/19 at 1000
	Nice
	Monaco for 1 night
	Menton for 1 night
	Imperia for 1 night
	Calvi for 1 night
	Propriano for 1 night
	Banifacio for 1 night
	Gallura for 1 night
	Maddalena for 1 night
	Cervo for 1 night
	Arbatax for 1 night
	Cagliari for 1 night
	Capri for 1 night
	Naples for 1 night
	crew wp leaves on 2/6/19 in Naples
	crew rb leaves on 2/6/19 in Naples


cruise  "Naples to Genoa via Amalfi Coast and Cinque Terre" departs Naples on 4/6/19 at 1000
	crew kmt joins on 2/6/19 in Naples
	crew sgr joins on 2/6/19 in Naples
	Naples
	Sorrento for 1 night
	Termini for 1 night
	Amalfi for 1 night
	Salerno for 1 night
	Capri for 1 night
	Ischia for 1 night
	Formia for 1 night
	Anzio for 1 night
	Ostia for 1 night
	Fanciullo for 1 night
	Orbetello for 1 night
	Follonica for 1 night
	Piombino for 1 night
	Portoferraio for 1 night
	Livorno for 1 night
	La_Spezia for 1 night
	Chiavari for 1 night
	Genoa
	crew smr leaves on 30/6/19 in Genoa
	crew isf leaves on 30/6/19 in Genoa
	crew po leaves on 30/6/19 in Genoa
	crew kmt leaves on 30/6/19 in Genoa
	crew sgr leaves on 30/6/19 in Genoa
