location IV_1 at 5 44'.37E 43 4'.66N is "W of Seche de Magnons Embiez"
location IV_2 at 5 51'.56E 43 2'.24N is "S of Cap Sicie"
location IV_3 at 5 57'.47E 43 4'.13N is "E of Cap Cepet light"
location IV_4 at 6 9'.14E 43 0'.68N is "Mid-channel Petite Passe"
location IV_5 at 6 12'.4E 42 58'.0N is "S of Cap dArmes"
location IV_6 at 6 21'.8E 43 4'.3N is "S of Cap Blanc Lighthouse"
location IV_7 at 6 33'.8E 43 3'.0N is "E of LeTitan"
