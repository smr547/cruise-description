vessel Trilogy name: "Trilogy" flag: "Australia" rego: 12345

location Sant_Carles is "Sant Carles de la Rapita"
location Barcelona is "Port of Barcelona Spain"
location Tarragona is "Port of Tarragona Spain"
location Blanes is "Blanes Spain"
location WPa at 6.7 43.2 is "a waypoint"
location Roses is "Roses Spain"
location Menton is "Menton Italy"
location Nice is "Port de Villefranche-sur-Mer, France"
location Cerbre is "Cape Cerbre France"
location Toulon is "Toulon France"
location Hyeres is "Hyeres France"
location Frejus is "Frejus France"
location Cannes is "Cannes France"
location Vendres is "Port Vendres"
location Bastia is "Bastia Corsica"
location Calvi is "Calvi Corsica"
location Macinaggio is "Macinaggio Corsica"
location Propriano is "Propriano Corsica"
location Banifacio is "Banifacio Corsica"
location Porto_Vecchio is "Porto Vecchio Corsica"
location ST_FLOR is "St Florent Corsica"
location Alghero is "Alghero Sardinia"
location Arbatax is "Arbatax Sardinia"
location Cagliari is "Cagliari Sardinia"
location Calsetta is "Calasetta Sardinia"
location Carloforte is "Carloforte Sardinia"
location Castelsardo is "Castelsardo Sardina"
location Rossa is "Isola Rossa Sardina"
location Maddalena is "Maddalena Archipelago Sardina"
location Olbia is "Olbia Sardinia"
location Cervo is "Porto Cervo Sardinia"
location Torres is "Porto Torres Sardinia"
location Portoscuso is "Portoscuso Sardinia"
location Gallura is "Santa Teresa Gallura Sardinia"
location Torregrande is "Torregrande  Sardinia"
location Tuelada is "Tuelada Sardinia"
location Villasimius is "Villasimius Sardinia"
location Imperia is "Imperia Italy"
location La_Spezia is "La Spezia Italy"
location Fanciullo is "Fanciullo Italy"
location Naples is "Naples Italy"
location Sorrento is "Sorrento Italy"
location Termini is "Termini Italy"
location Amalfi is "Amalfi Italy"
location Salerno is "Salerno Italy"
location Capri is "Capri Italy"
location Ischia is "Ischia Italy"
location Formia is "Formia Italy"
location Anzio is "Anzio Italy"
location Ostia is "Ostia Italy"
location Orbetello is "Orbetello Italy"
location Follonica is "Follonica Italy"
location Piombino is "Piombino Italy"
location Portoferraio is "Portoferraio Italy"
location Livorno is "Livorno Italy"
location Chiavari is "Chiavari Italy"
location Genoa is "Genoa Italy"
location Monaco is "Monaco"

person smr name: "Steven Michael Ring"
person isf name: "Irene Sarah Farthing"
person po name: "Peter Olaf Otteson"
person gh name: "Graeme Hubbard"
person sm name: "Cheryl Meikle"
person sjr name: "Steven James Ring"
person pjr name: "Patrick James Ring"
person ar name: "Alice Ring"
person kmt name: "Karyn Marie Talty"
person sgr name: "Stephen Gordon Reeves"
person wp name: "Wayne Petschack"
person rb name: "Rena Brettle"

season Steven_cruise vessel Trilogy begins in Sant_Carles

cruise  "Shakedown" departs Sant_Carles on 14/4/19
	Sant_Carles
        crew smr joins on 31/3/19 as skipper in Sant_Carles
        crew wp  joins on 08/4/19 as mate in Sant_Carles
	Tarragona for 1 night
	Barcelona for 4 nights
        crew wp leaves on 16/4/19

cruise  "Barcelona to Nice" departs Barcelona on 14/4/19
        crew gh joins on 16/4/19 in Barcelona
        crew cm joins on 16/4/19 in Barcelona
        crew sjr joins on 16/4/19 in Barcelona
        crew pjr joins on 16/4/19 in Barcelona
        crew ar joins on 16/4/19 in Barcelona
	Barcelona
	Blanes for 1 night
	Roses for 1 night
	Cerbre for 1 night
	Vendres for 1 night
	Toulon for 1 night
	Hyeres for 1 night
	WPa
	Frejus for 1 night
	Cannes for 1 night
	Nice for 4 nights
	crew gh leaves on 30/4/19 in Nice
	crew cm leaves on 30/4/19 in Nice
	crew sjr leaves on 1/5/19 in Nice
	crew ar leaves on 1/5/19 in Nice
	crew pjr leaves on 1/5/19 in Nice

cruise  "Nice to Naples via Corsica and Sardinia" departs Nice on 3/5/19
	crew po joins on 1/5/19 as mate in Nice
	crew wp joins on 1/5/19 in Nice
	crew rb joins on 1/5/19 in Nice
	crew isf joins on 2/5/19 in Nice 
	Nice
	Monaco for 1 night
	Menton for 1 night
	Imperia for 1 night
	Calvi for 1 night
	Propriano for 1 night
	Banifacio for 1 night
	Gallura for 1 night
	Maddalena for 1 night
	Cervo for 1 night
	Arbatax for 1 night
	Cagliari for 1 night
	Capri for 1 night
	Naples for 1 night
	crew wp leaves on 2/6/19 in Naples
	crew rb leaves on 2/6/19 in Naples


cruise  "Naples to Genoa via Amalfi Coast and Cinque Terre" departs Naples on 4/6/19
	crew kmt joins on 2/6/19 in Naples
	crew sgr joins on 2/6/19 in Naples
	Naples
	Sorrento for 1 night
	Termini for 1 night
	Amalfi for 1 night
	Salerno for 1 night
	Capri for 1 night
	Ischia for 1 night
	Formia for 1 night
	Anzio for 1 night
	Ostia for 1 night
	Fanciullo for 1 night
	Orbetello for 1 night
	Follonica for 1 night
	Piombino for 1 night
	Portoferraio for 1 night
	Livorno for 1 night
	La_Spezia for 1 night
	Chiavari for 1 night
	Genoa
	crew smr leaves on 30/6/19 in Genoa
	crew isf leaves on 30/6/19 in Genoa
	crew po leaves on 30/6/19 in Genoa
	crew kmt leaves on 30/6/19 in Genoa
	crew sgr leaves on 30/6/19 in Genoa
