person smr name: "Steven Michael Ring"
person isf name: "Irene Sarah Farthing"
person po name: "Peter Olaf Otteson"
person gh name: "Graeme Hubbard"
person cm name: "Cheryl Meikle"
person sjr name: "Steven James Ring"
person pjr name: "Patrick James Ring"
person ar name: "Alice Ring"
person kmt name: "Karyn Marie Talty"
person sgr name: "Stephen Gordon Reeves"
person wp name: "Wayne Petschack"
person rb name: "Rena Brettle"
person eif name: "Emily Farthing"
person pl name: "Peter Lucey"
person sl name: "Sue Lucey"
person tt name: "Theo Theodosi"
person lt name: "Lana Theodosi"
