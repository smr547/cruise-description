vessel Trilogy name: "Trilogy" flag: "Australia" rego: 12345 speed: 7.5

use http://planacruise.online/locations/spain_med_coast.txt
use http://planacruise.online/locations/sardinia.txt
use http://planacruise.online/locations/sicily.txt
use http://planacruise.online/locations/balearics.txt
use http://planacruise.online/locations/north_africa.txt
use http://planacruise.online/locations/malta.txt

use file:///Users/stevenring/projects/cruise-description/grammar/people.cdl

season steven_2020 vessel Trilogy begins in Sant_Carles

# smr and isf arrive Barcelona Monday 23 March at 6:30am then bus to Sant Carles arriving around Midday
# smr will conduct hull inspections to ensure antifoul, anodes, saildrive foot and other preparations are satisfactory prior to relaunch
# if all is satisfactory, Trilogy will be relaunch on 24 March 2020 at Sant Carles Marina


cruise  "Shakedown - Sant Carles to Tarragona" departs Sant_Carles on 2/4/20 at 1000
	Sant_Carles
        crew smr joins on 23/3/20 as skipper in Sant_Carles
        crew isf joins on 23/3/20 in Sant_Carles
        crew wp joins on 25/3/20 as mate in Sant_Carles
	via Calafat
        Tarragona for 1 night

cruise  "Passage - Tarragona to Majorca" departs Tarragona on 3/4/20 at 1600
	Tarragona
        Soller for 3 nights


cruise  "Cruising Majorca" departs Soller on 7/4/20 at 1000
        Soller
	via Sant_Elm
	Camp_de_Mar for 1 night
	via Sol_de_Mallorca
        Palma for 2 nights
	Cabrera for 1 night
	via Cala_Millor
        Alcudia for 1 night


cruise  "Cruising Menorca" departs Alcudia on 12/4/20 at 0800
	Alcudia
	Ciutadella for 1 night
	via Xoriguer
	Serpentona for 1 night
	via Punta_Prima
        Mahon for 2 nights

cruise  "Passage - Menorca to Sardina" departs Mahon on 17/4/20 at 0900
	Mahon
	Alghero for 2 nights
        crew rb joins on 18/4/20 in Alghero

cruise  "Cruising Sardina" departs Alghero on 19/4/20 at 0800
	Alghero
	Bosa for 1 night
	Torregrande for 2 nights 
        Portoscuso for 1 night
        Carloforte for 1 night
        Calsetta for 1 night
        Tuelada for 1 night
	Cagliari for 3 night
        crew rb leaves

cruise  "Passage - Sardina to Tunisia" departs Cagliari on 27/4/20 at 1000
        Cagliari
        Goulette for 3 nights


cruise  "Passage - Tunisa to Silicy" departs Goulette on 1/5/20 at 1300
	Goulette
        Marsala for 3 nights
        crew rb joins on 2/5/20 in Marsala

cruise "North Sicily" departs Marsala on 5/5/20 at 1000
	Marsala
	Trapani for 2 nights
        Palermo for 3 nights
        Cefalu for 2 nights
        Gregorio for 3 nights

cruise "Aeolian Islands" departs Gregorio on 15/5/20 at 0900
	Gregorio
	Lipari for 12 nights
        crew wp leaves
        crew rb leaves


cruise "South Sicily" departs Lipari on 26/5/20 at 1000
	Lipari
        Messina for 3 nights
        Catania for 3 nights
        Siracusa for 3 nights
	Pozzallo for 3 nights
	Gela for 3 nights
        Licata for 2 nights
        Empedocle for 2 nights

cruise "Sicily to Malta" departs Empedocle on 17/6/20 at 1700
	Empedocle
	Marsalforn for 1 night

cruise "Malta Miandering" departs Marsalforn on 19/6/20 at 1000
	Marsalforn
	Mgarr for 1 night
	Blue_Lagoon for 1 night
	Santa_Marija for 1 night
	Mellieha for 1 night
	Portomaso for 1 nights
	Valetta for 3 nights
        crew smr leaves
        crew isf leaves
